// ��λ, �����һ����λ���ֺ�һ����λ���ְ�λ�߼�����, ��Ҫ����λ����replacateΪ��λ���ֵĳ���
// e.g. b[15:0]^{16{sub}}

// ->(H)casez, casex: z��x������Ϊͨ���ʹ��
// concentration  previlege

// ->(H) ��ǰ��Ĭ��ֵ

// ->(H) ��������ʵ��  generate + for 
/*
module top_module( 
    input [99:0] a, b,
    input cin,
    output [99:0] cout,
    output [99:0] sum );
    

    full_adder adder0(.cin(cin), .cout(cout[0]), .a(a[0]), .b(b[0]), .sum(sum[0]));
    genvar i;
    generate 
        for(i = 1; i < 100; i++) begin: all_adder
            full_adder adder(.cin(cout[i-1]), .cout(cout[i]), .a(a[i]), .b(b[i]), .sum(sum[i]));           
        end
    endgenerate
                             
            
endmodule
*/

// ->(H) reg�Ĵ����޷�ֱ�Ӹ���ʼֵ, ֻ���ڵ�һ��ʱ��(�ϵ�)��ʱ����һ��reset�ź���always�������� 

// ->(H) {pm, hh, mm, ss} = {1'b0, 8'd12, 8'd0, 8'd0}
//       �����ַ�����ֵʱ, ����Ҫд���λ��
//       ����ʱ��Ҳһ��, λ����ʽ��

// ->(H) ʵ�� �в㼶��������˳���״̬ת��
//       if, case, ?:�����϶�������, ���Ǻ�����ֻ���ǲ���,
//       for������ʱ�Ӳ�����, ����Ƕ��ֻ����if
        /*
        ��һ�� always @(posedge clk) ��ʱ����
        ���Ҫ���в㼶��������˳���״̬ת�ƣ�Ƕ���㷨������
        ʵ����ֻ���� if / else Ƕ�ס�
        */

