
// ���� ��дverilog��ʱ��, ע�� ǿĿ��������, �γɷ��, �γ�ϰ��    ���ռ�����ʦ��Ҫ��
//    -------����ע�⼸��--------
/*
1. �����߼���·����
2. ��Ӧ�߼���·���ص�, ǿĿ����������ѡ�����Ƶ�д��, �����γ���Ʒ���ϰ��

*/

/*
1---> Key Words:
module
input output
assign always
endmodule
*/

/*
2---> Basic Operators in Verilog (bitwise/logical/reduction/case):
~      bitwise NOT
!      logical NOT

& | ^        bitwise AND OR XOR
&& ||        logical AND OR

~& ~| ~^     bitwise NAND NOR XNOR

&a |a ^a     reduction AND OR XOR
~&a ~|a ~^a  reduction NAND NOR XNOR

== !=        logical equality
=== !==      case equality

others:
{}      concatenation
{}:n    replication
?:      conditional
*/


/*
3---> Variables in Verilog:
wire                       represents physical connections
reg                        represents storage elements (flip-flops) ��:ֻ����always�����渳ֵ
integer                    ���ڸ�������������, ��ѭ��i

vector [m:n]               represents multiple bits (m>n)
*/

/*
4 ---> Number representaion:
N'bXXXX      N bits binary
N'dXXXX      N bits decimal
N'hXXXX      N bits hexadecimal
N'oXXXX      N bits octal
*/

/*
5 ---> functions::
if   case  for    generate + for
*/

/*
6 ---> System function:
$bits(variable)          returns the size (in bits) of the variable
*/


/*
7 ---> Write Testbench:
testbench���Խű�����Ӳ��, ֻ�ǽű�, initial���о��ǽű�����
`timescale ../..
initial forever

����ʱ��:
`timescale 1ps/1ps
module top_module ( );
    reg clk;

    // 1?? ʵ���� DUT��ʵ�������⣬������ u_dut��
    dut u_dut (
        .clk(clk)
        // �����˿�����У������Ȳ�������
    );

    // 2?? ʱ�Ӳ��������� 10 ps����ʼΪ 0����һ��������
    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;  // 5 ps ��תһ�� �� ���� 10 ps
    end
endmodule

���첨��:
module top_module ( output reg A, output reg B );//

    // generate input patterns here
    initial begin
        A = 0; B = 0;
        #10 A = 1;
        #5  B = 1;
        #5 A = 0;
        #20 B = 0;
    end


endmodule

`timescale 1ps/1ps
module top_module();
    reg clk;
    reg in;
    reg [2:0] s;
    wire out;
    
    q7 test_q7(.clk(clk), .in(in), .s(s), .out(out));
    
    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        in = 1'b0;
        s = 3'b010;
        #10 s = 3'b110;
        #10 begin
            s = 3'b010;
            in = 1;
        end
        #10 begin
            s = 3'b111;
            in = 0;
        end
        #10 begin
            s = 3'b000;
            in = 1;
        end
        #30 in = 0;
    end

endmodule
*/