// module-module name-input&output   endmodule   
/*
module-moduleName-(�˿��б�);
�˿��ź����� (�����������, �źŵ���������, �źŵ�λ��); 
input output inout; wire reg logic; λ��[n1:n2]
�������� parameter ...
*/
// assign �ڲ��ź�����

// always �ײ�ģ�����ԭ�����
/*
@ means "at", "wait for", ��ֵ���� must be reg type     (begin end ֮����˳��ִ��, ������ִ��)
negedge posedge �½���, ������      
e.g. always @(D);  // whenever D changes excute the command
��: if case for , could be used in always block
һ����˵ʱ���߼���ֵҪ�� A <= B;  // non-blocking assignment  ��������ֵ
����߼���ֵҪ�� A = B;   // blocking assignment  ������ֵ
��:һ�� always ����ֻ����һ�ָ�ֵ��ʽ
*/

// ��ԭ��: ���� and or xor ... ����ֱ����, �����Ͼ����Ѿ���װ�õĵײ�ģ��

// ��������:
// net�е���������: wire tri supply0....                     ��wireΪ��
// variable�е���������: reg integer time real realtime...   ��regΪ��

// ���ֱ�ʾ:
// 6' b010100    8' sb10010111 = -010111   5' d14 = 01110 

// �߼�(bool)��ʾ:
// 1, 0, x, z(����̬)

//-------------------------------
// ����verilog������:
// �ŵ�·��: ֱ������, ���ǹ��ڷ�װ, ���Ժ��ײ��߼�, д���������ֱ�ӻ�ԭ��ͼ. ���ȼ�(3)
// assign��: ��������֮��, һ���Ǵ�����߼�ʵ�������, д��������������߼�����. ���ȼ�(2)
// always��: �ȽϺõ�һ�����ֱ�ӿ�����if case for, �����߼��Ѻ�. ���ȼ�(1)

// module structure test:
module MUX2to1(
    input wire A, 
    input wire B,
    input wire Sel,
    output wire Y
)
assign Y = Sel ? B : A;
endmodule

module edge_DFF(
    input wire D,
    input wire CLK,
    output reg Q,
    output reg Qbar
)
always @(posedge CLK)   
begin
    Q <= D;
    Qbar <= ~D;
end
endmodule

module full_subtractor();

endmodule

module random_test(A, B, Y);
    input wire A;
    input wire B;
    output wire Y;

    assign M = A !&& B;
    assign T = A ~^ M;
    assign Y = T !|| B;
endmodule 

module full_adder(A, B, Carry_in, S, Carry_out);
    input wire [3:0] A, B;
    input wire Carry_in;
    output reg [3:0] S;
    output reg Carry_out;

endmodule


// logic words test:

Y = ~8' b10101000;






