
// ���� ��дverilog��ʱ��, ע�� ǿĿ��������, �γɷ��, �γ�ϰ��    ���ռ�����ʦ��Ҫ��
//    -------����ע�⼸��--------
/*
1. �����߼���·����
2. ��Ӧ�߼���·���ص�, ǿĿ����������ѡ�����Ƶ�д��, �����γ���Ʒ���ϰ��

*/

/*
1---> Key Words:
module
input output
assign always
endmodule
*/

/*
2---> Basic Operators in Verilog (bitwise/logical/reduction/case):
~      bitwise NOT
!      logical NOT

& | ^        bitwise AND OR XOR
&& ||        logical AND OR

~& ~| ~^     bitwise NAND NOR XNOR

&a |a ^a     reduction AND OR XOR
~&a ~|a ~^a  reduction NAND NOR XNOR

== !=        logical equality
=== !==      case equality

others:
{}      concatenation
{}:n    replication
?:      conditional
*/


/*
3---> Variables in Verilog:
wire                       represents physical connections
reg                        represents storage elements (flip-flops) ��:ֻ����always�����渳ֵ
integer                    ���ڸ�������������, ��ѭ��i

vector [m:n]               represents multiple bits (m>n)
*/

/*
4 ---> Number representaion:
N'bXXXX      N bits binary
N'dXXXX      N bits decimal
N'hXXXX      N bits hexadecimal
N'oXXXX      N bits octal
*/

/*
5 ---> functions::
if   case  for    generate + for
*/

/*
6 ---> System function:
$bits(variable)          returns the size (in bits) of the variable
*/
