// ��λ, �����һ����λ���ֺ�һ����λ���ְ�λ�߼�����, ��Ҫ����λ����replacateΪ��λ���ֵĳ���
// e.g. b[15:0]^{16{sub}}

// ->(H)casez, casex: z��x������Ϊͨ���ʹ��
// concentration  previlege

// ->(H) ��ǰ��Ĭ��ֵ

// ->(H) ��������ʵ��  generate + for 
/*
module top_module( 
    input [99:0] a, b,
    input cin,
    output [99:0] cout,
    output [99:0] sum );
    

    full_adder adder0(.cin(cin), .cout(cout[0]), .a(a[0]), .b(b[0]), .sum(sum[0]));
    genvar i;
    generate 
        for(i = 1; i < 100; i++) begin: all_adder
            full_adder adder(.cin(cout[i-1]), .cout(cout[i]), .a(a[i]), .b(b[i]), .sum(sum[i]));           
        end
    endgenerate
                             
            
endmodule
*/

// ->(H) reg�Ĵ����޷�ֱ�Ӹ���ʼֵ, ֻ���ڵ�һ��ʱ��(�ϵ�)��ʱ����һ��reset�ź���always�������� 

// ->(H) {pm, hh, mm, ss} = {1'b0, 8'd12, 8'd0, 8'd0}
//       �����ַ�����ֵʱ, ����Ҫд���λ��
//       ����ʱ��Ҳһ��, λ����ʽ��

// ->(H) ʵ�� �в㼶��������˳���״̬ת��
//       if, case, ?:�����϶�������, ���Ǻ�����ֻ���ǲ���,
//       for������ʱ�Ӳ�����, ����Ƕ��ֻ����if
        /*
        ��һ�� always @(posedge clk) ��ʱ����
        ���Ҫ���в㼶��������˳���״̬ת�ƣ�Ƕ���㷨������
        ʵ����ֻ���� if / else Ƕ�ס�
        */

// ->   ��Ϊ if  elseif elseif... else����һ�ױ��������Ⱥ��ϵ, ���Կ��Բ���ififif...Ƕ��

// ->   ʹ�� one-hot ״̬�����������: ����FSM��ʵ��, ���Ը������ʹ�ù�ȥ�Ƶ���״̬, 
//      һ����˵״̬����ֱ�۵ط����϶�����������next_state
// e.g.
/*
module top_module(
    input in,
    input [3:0] state,
    output [3:0] next_state,
    output out); //

    parameter A=0, B=1, C=2, D=3;

    // State transition logic: Derive an equation for each state flip-flop.
    assign next_state[A] = state[A] & ~in | state[C] & ~in;
    assign next_state[B] = state[A] & in | state[B] & in | state[D] & in;
    assign next_state[C] = state[B] & ~in | state[D] & ~in;
    assign next_state[D] = state[C] & in;

    // Output logic: 
    assign out = (state[D] == 1);

endmodule
*/

// ->(H)
/*
FSM�Ŀ����������Ҫ�ֶ�����, ��ô���������state���и���, �����Գ�״̬. 
��״̬ѭ��������, ���ʱ�ѿ����������Ϳɸ�ԭ�Ժ�������
���������¾��Բ���������, ����״̬����, ������������״̬��

reset��Ҫע��ʵʱ��, ����Ӧ������Ϊһ��ʱ���������ʱһ��ʱ����Ч, ����Ҫ������жϼ�ʱ��Ч
*/

// ->(H) ����Ǵ��ܽ�, ���Զ��������ϵͳ�����������:
/*
ϵͳ���ʱ�ķֿ�����:
��Ϻ�datapath������÷ֿ�
ʱ�򲿷�: ���Բ��д��зֿ�, 
������ˮ�߷ֿ��ǹ��̱�׼��(����һ�����������Ϊ��һ���Ŀ�����)
Ƕ�׷ֿ��ʱ��Ҫע������ʱ��

���ĵײ�ģ��ֻ��������, ��д�߼�, ����������ά��.
*/

// ���м��ģ��
// module seq_1101 (
//     input  clk,
//     input  reset,
//     input  data,
//     output start
// );

//     typedef enum logic [2:0] {
//         S0, S1, S11, S110
//     } state_t;

//     state_t state, next;

//     always @(posedge clk) begin
//         if (reset)
//             state <= S0;
//         else
//             state <= next;
//     end

//     always @(*) begin
//         case (state)
//             S0:   next = data ? S1   : S0;
//             S1:   next = data ? S11  : S0;
//             S11:  next = data ? S11  : S110;
//             S110: next = data ? S1   : S0;   // overlap ok
//             default: next = S0;
//         endcase
//     end

//     // Mealy pulse on detecting 1101
//     assign start = (state == S110) && data;

// endmodule


// module timer_fsm (
//     input  clk,
//     input  reset,
//     input  start,
//     input  done_counting,
//     input  ack,
//     output shift_ena,
//     output counting,
//     output done
// );

//     typedef enum logic [1:0] {
//         RECOG,
//         SHIFT,
//         COUNT,
//         DONE
//     } state_t;

//     state_t state, next;

//     // shift counter (FSM-owned)
//     reg [1:0] shift_cnt;

//     // state + counter register
//     always @(posedge clk) begin
//         if (reset) begin
//             state     <= RECOG;
//             shift_cnt <= 2'd0;
//         end else begin
//             state <= next;

//             if (state == SHIFT)
//                 shift_cnt <= shift_cnt + 1'b1;
//             else
//                 shift_cnt <= 2'd0;
//         end
//     end

//     // next-state logic
//     always @(*) begin
//         case (state)
//             RECOG: next = start ? SHIFT : RECOG;

//             SHIFT: next = (shift_cnt == 2'd3) ? COUNT : SHIFT;

//             COUNT: next = done_counting ? DONE : COUNT;

//             DONE:  next = ack ? RECOG : DONE;

//             default: next = RECOG;
//         endcase
//     end

//     // outputs (pure Moore)
//     assign shift_ena = (state == SHIFT);
//     assign counting  = (state == COUNT);
//     assign done      = (state == DONE);

// endmodule


// // ����ģ��ֻ����, ��ģ�鶼д��, ����ֻ��ģ��.  �����hierarchyҲһ��, ÿһ��ģ��Ķ��㶼��ֻ����, ��ʵ���߼�
// module top_module (
//     input  clk,
//     input  reset,
//     input  data,
//     output shift_ena,
//     output counting,
//     input  done_counting,
//     output done,
//     input  ack
// );

//     wire start;
//     wire seq_recog_reset;

//     seq_1101 u_seq (
//         .clk   (clk),
//         .reset(reset),
//         .data  (data),
//         .start (start)
//     );

//     timer_fsm u_fsm (
//         .clk          (clk),
//         .reset        (reset),
//         .start        (start),
//         .done_counting(done_counting),
//         .ack          (ack),
//         .shift_ena    (shift_ena),
//         .counting     (counting),
//         .done         (done)
//     );

// endmodule

